class seq;
endclass
