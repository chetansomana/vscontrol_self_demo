class gpio_seq;

  input bit a;
  output bit b;
endclass
