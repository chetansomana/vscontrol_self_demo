class
class
class
class
