class
class
